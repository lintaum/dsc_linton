`define ADDR_WIDTH 7
`define FONTE 32'd0
`define DESTINO 32'd75
`define CUSTO_CAMINHO 32'd47
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd11
`define MAX_ATIVOS 32'd13
`define TAMANHO_CAMINHO 13
`define MENOR_CAMINHO {7'd0, 7'd1, 7'd10, 7'd18, 7'd17, 7'd24, 7'd32, 7'd41, 7'd49, 7'd57, 7'd65, 7'd74, 7'd75}