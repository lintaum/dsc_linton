`define ADDR_WIDTH 6
`define FONTE 32'd0
`define DESTINO 32'd41
`define CUSTO_CAMINHO 32'd38
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd10
`define MAX_ATIVOS 32'd9
`define TAMANHO_CAMINHO 12
`define MENOR_CAMINHO {6'd0, 6'd1, 6'd8, 6'd14, 6'd13, 6'd20, 6'd25, 6'd31, 6'd32, 6'd27, 6'd34, 6'd41}