`define ADDR_WIDTH 6
`define FONTE 32'd0
`define DESTINO 32'd37
`define CUSTO_CAMINHO 32'd32
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd10
`define MAX_ATIVOS 32'd9
`define TAMANHO_CAMINHO 9
`define MENOR_CAMINHO {6'd0, 6'd1, 6'd8, 6'd14, 6'd13, 6'd20, 6'd25, 6'd30, 6'd37}