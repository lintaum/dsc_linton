`define ADDR_WIDTH 7
`define FONTE 32'd0
`define DESTINO 32'd111
`define CUSTO_CAMINHO 32'd57
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd11
`define MAX_ATIVOS 32'd19
`define TAMANHO_CAMINHO 13
`define MENOR_CAMINHO {7'd0, 7'd1, 7'd11, 7'd22, 7'd32, 7'd41, 7'd52, 7'd61, 7'd71, 7'd80, 7'd90, 7'd100, 7'd111}