`define ADDR_WIDTH 10
`define FONTE 10'd0
`define DESTINO 10'd98
`define CUSTO_CAMINHO 10'd54
`define MAX_ATIVOS 10'd17
`define TAMANHO_CAMINHO 12
`define MENOR_CAMINHO {10'd0, 10'd1, 10'd11, 10'd21, 10'd30, 10'd40, 10'd49, 10'd59, 10'd69, 10'd79, 10'd88, 10'd98}