`define ADDR_WIDTH 10
`define FONTE 32'd0
`define DESTINO 32'd1022
`define CUSTO_CAMINHO 32'd179
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd14
`define MAX_ATIVOS 32'd61
`define TAMANHO_CAMINHO 60
`define MENOR_CAMINHO {10'd0, 10'd31, 10'd63, 10'd95, 10'd127, 10'd159, 10'd160, 10'd192, 10'd193, 10'd163, 10'd164, 10'd165, 10'd166, 10'd167, 10'd198, 10'd230, 10'd200, 10'd201, 10'd233, 10'd265, 10'd266, 10'd235, 10'd205, 10'd206, 10'd238, 10'd269, 10'd301, 10'd333, 10'd365, 10'd396, 10'd427, 10'd458, 10'd490, 10'd521, 10'd552, 10'd583, 10'd615, 10'd645, 10'd676, 10'd707, 10'd706, 10'd736, 10'd766, 10'd798, 10'd829, 10'd859, 10'd827, 10'd857, 10'd888, 10'd920, 10'd952, 10'd984, 10'd1015, 10'd985, 10'd986, 10'd1018, 10'd1019, 10'd989, 10'd1021, 10'd1022}