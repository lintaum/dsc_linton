`define ADDR_WIDTH 7
`define FONTE 32'd0
`define DESTINO 32'd69
`define CUSTO_CAMINHO 32'd53
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd11
`define MAX_ATIVOS 32'd15
`define TAMANHO_CAMINHO 10
`define MENOR_CAMINHO {32'd0, 32'd8, 32'd16, 32'd25, 32'd26, 32'd35, 32'd43, 32'd52, 32'd60, 32'd69}