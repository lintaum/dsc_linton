`define ADDR_WIDTH 4
`define FONTE 32'd0
`define DESTINO 32'd14
`define CUSTO_CAMINHO 32'd24
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd8
`define MAX_ATIVOS 32'd3
`define TAMANHO_CAMINHO 5
`define MENOR_CAMINHO {4'd0, 4'd3, 4'd7, 4'd11, 4'd14}