`define ADDR_WIDTH 10
`define FONTE 32'd0
`define DESTINO 32'd1021
`define CUSTO_CAMINHO 32'd158
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd14
`define MAX_ATIVOS 32'd64
`define TAMANHO_CAMINHO 60
`define MENOR_CAMINHO {10'd0, 10'd1, 10'd33, 10'd64, 10'd96, 10'd66, 10'd67, 10'd98, 10'd130, 10'd162, 10'd194, 10'd164, 10'd165, 10'd166, 10'd136, 10'd137, 10'd169, 10'd200, 10'd201, 10'd233, 10'd265, 10'd266, 10'd267, 10'd299, 10'd331, 10'd332, 10'd302, 10'd303, 10'd335, 10'd365, 10'd395, 10'd425, 10'd455, 10'd486, 10'd518, 10'd550, 10'd582, 10'd613, 10'd643, 10'd675, 10'd705, 10'd737, 10'd768, 10'd798, 10'd829, 10'd828, 10'd827, 10'd857, 10'd888, 10'd920, 10'd952, 10'd984, 10'd1015, 10'd985, 10'd986, 10'd1018, 10'd1019, 10'd1020, 10'd989, 10'd1021}