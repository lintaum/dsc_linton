`define ADDR_WIDTH 11
`define FONTE 32'd0
`define DESTINO 32'd2046
`define CUSTO_CAMINHO 32'd208
`define CUSTO_WIDTH 32'd4
`define MAX_VIZINHOS 32'd8
`define DISTANCIA_WIDTH 32'd15
`define MAX_ATIVOS 32'd80
`define TAMANHO_CAMINHO 54
`define MENOR_CAMINHO {11'd0, 11'd1, 11'd47, 11'd93, 11'd138, 11'd183, 11'd227, 11'd272, 11'd318, 11'd319, 11'd365, 11'd410, 11'd456, 11'd502, 11'd547, 11'd591, 11'd635, 11'd679, 11'd725, 11'd770, 11'd816, 11'd862, 11'd908, 11'd953, 11'd952, 11'd996, 11'd1042, 11'd1088, 11'd1134, 11'd1180, 11'd1181, 11'd1227, 11'd1271, 11'd1316, 11'd1361, 11'd1407, 11'd1453, 11'd1498, 11'd1544, 11'd1589, 11'd1633, 11'd1678, 11'd1679, 11'd1725, 11'd1726, 11'd1772, 11'd1818, 11'd1864, 11'd1863, 11'd1908, 11'd1954, 11'd1999, 11'd2045, 11'd2046}